module Top_Module_tb;

    timeunit 1ns/1ps;

    logic SC_EN = 0;
    logic clk   = 0;

   
    logic [15:0] pgm [0:255];


    logic prog_wr_en;
    logic [11:0] prog_addr;
    logic [15:0] prog_data;
  	logic rst;
  logic [7:0] input_data;
  logic input_read;
  logic [11:0]PC_Reset_Initial_Data;
  	logic PC_Reset_Initial;

    Top_Module CPU (
        .clk(clk),
        .SC_EN(SC_EN),
      	.rst(rst),
        .prog_wr_en(prog_wr_en),
        .prog_addr(prog_addr),
      .prog_data(prog_data),
      .input_data(input_data),
      .input_read(input_read),
      .PC_Reset_Initial_Data(PC_Reset_Initial_Data),
      .PC_Reset_Initial(PC_Reset_Initial)      
    );

    localparam clk_period = 10;

    
    initial begin
        forever begin
          #(clk_period/2) clk = ~clk;
          
        end
    end

    
    initial begin
      PC_Reset_Initial_Data = 12'b0;
      pgm[0]  = 16'h7800;
      pgm[1]  = 16'h504F;
      pgm[2]  = 16'h3014;
      pgm[3]  = 16'h2012;
      pgm[4]  = 16'h7200;
      pgm[5]  = 16'h7020;
      pgm[6]  = 16'h1014;
      pgm[7]  = 16'h7004;
      pgm[8]  = 16'h400A;
      pgm[9]  = 16'h4016;
      pgm[10]  = 16'h5022;
      pgm[11]  = 16'h3013;
      pgm[12]  = 16'h2021;
      pgm[13]  = 16'h7800;
      pgm[14]  = 16'h3021;
      pgm[15]  = 16'h5034;
      pgm[16]  = 16'hB013;
      pgm[17]  = 16'h4000;
      pgm[18]  = 16'h0010;
      pgm[19]  = 16'h0000;
      pgm[20]  = 16'h0000;
      pgm[21]  = 16'h0000;
      pgm[22]  = 16'h5034;
      pgm[23]  = 16'h3015;
      pgm[24]  = 16'hC015;
      pgm[25]  = 16'hfff0;
      pgm[26]  = 16'h0000;
      pgm[27]  = 16'h7040;
      pgm[28]  = 16'h7040;
      pgm[29]  = 16'h7040;
      pgm[30]  = 16'h7040;
      pgm[31]  = 16'h0019;
      pgm[32]  = 16'hC01A;
      pgm[33]  = 16'h0000;
      pgm[34]  = 16'h0000;
      pgm[35]  = 16'h2014;
      pgm[36]  = 16'h501A;
      pgm[37]  = 16'h3021;
      pgm[38]  = 16'h7800;
      pgm[39]  = 16'h504F;
      pgm[40]  = 16'h1021;
      pgm[41]  = 16'h501A;
      pgm[42]  = 16'h3021;
      pgm[43]  = 16'h7800;
      pgm[44]  = 16'h504F;
      pgm[45]  = 16'h1021;
      pgm[46]  = 16'h501A;
      pgm[47]  = 16'h3021;
      pgm[48]  = 16'h7800;
      pgm[49]  = 16'h504F;
      pgm[50]  = 16'h1021;
      pgm[51]  = 16'hC022;
      pgm[52]  = 16'h0000;
      pgm[53]  = 16'h7800;
      pgm[54]  = 16'h504F;
      pgm[55]  = 16'h1021;
      pgm[56]  = 16'h501A;
      pgm[57]  = 16'h3021;
      pgm[58]  = 16'h7800;
      pgm[59]  = 16'h504F;
      pgm[60]  = 16'h1021;
      pgm[61]  = 16'h501A;
      pgm[62]  = 16'h3021;
      pgm[63]  = 16'h7800;
      pgm[64]  = 16'h504F;
      pgm[65]  = 16'h1021;
      pgm[66]  = 16'h501A;
      pgm[67]  = 16'h3021;
      pgm[68]  = 16'h7800;
      pgm[69]  = 16'h504F;
      pgm[70]  = 16'h1021;
      pgm[71]  = 16'hC034;
      pgm[72]  = 16'h0000;
      pgm[73]  = 16'h0039;
      pgm[74]  = 16'h0041;
      pgm[75]  = 16'h0030;
      pgm[76]  = 16'h000a;
      pgm[77]  = 16'h0020;
      pgm[78]  = 16'h000d;
      pgm[79]  = 16'h0000;
      pgm[80]  = 16'hF200;
      pgm[81]  = 16'h4050;
      pgm[82]  = 16'hF800;
      pgm[83]  = 16'h3048;
      pgm[84]  = 16'h204D;
      pgm[85]  = 16'h7200;
      pgm[86]  = 16'h7020;
      pgm[87]  = 16'h1048;
      pgm[88]  = 16'h7004;
      pgm[89]  = 16'h405B;
      pgm[90]  = 16'h4050;
      pgm[91]  = 16'h204E;
      pgm[92]  = 16'h7200;
      pgm[93]  = 16'h7020;
      pgm[94]  = 16'h1048;
      pgm[95]  = 16'h7004;
      pgm[96]  = 16'h4062;
      pgm[97]  = 16'h404F;
      pgm[98]  = 16'h2049;
      pgm[99]  = 16'h7200;
      pgm[100]  = 16'h7020;
      pgm[101]  = 16'h1048;
      pgm[102]  = 16'h7004;
      pgm[103]  = 16'h4069;
      pgm[104]  = 16'h4073;
      pgm[105]  = 16'h7040;
      pgm[106]  = 16'h7002;
      pgm[107]  = 16'h4073;
      pgm[108]  = 16'h406D;
      pgm[109]  = 16'h204A;
      pgm[110]  = 16'h7200;
      pgm[111]  = 16'h7020;
      pgm[112]  = 16'h1048;
      pgm[113]  = 16'h104C;
      pgm[114]  = 16'hC04F;
      pgm[115]  = 16'h204B;
      pgm[116]  = 16'h7200;
      pgm[117]  = 16'h7020;
      pgm[118]  = 16'h1048;
      pgm[119]  = 16'hC04F;
    end
  
  	integer i;

    
    initial begin
      	$dumpfile("dump.vcd"); $dumpvars(0, CPU);
      	input_read = 0;
      	rst = 1;
        SC_EN = 0;
        prog_wr_en = 0;
        prog_addr  = 0;
        prog_data  = 16'd0;
		#10
        @(posedge clk);
      	rst = 0;
      	PC_Reset_Initial = 1;
	
        
      for (i = 0; i < 120; i = i + 1) begin
            prog_wr_en = 1;
            prog_addr  = i;
            prog_data  = pgm[i];
            @(posedge clk);  
        end
      

        
      
      
            @(posedge clk);  
        
      	PC_Reset_Initial = 0;
        prog_wr_en = 0;
        SC_EN = 1;
        

        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "8";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "5";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "6";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "B";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "8";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "9";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "A";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "B";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "C";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "D";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "E";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "6";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "F";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "7";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "F";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "F";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "F";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "8";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "F";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "3";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "B";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "1";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "4";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h20;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'hD;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= 8'h47;
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "2";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;
        #2000 input_data <= "0";
        #1 input_read <= 1;
        #20 input_read <= 0;

      

        
      #20000 
      $display(" input buffer = %h", CPU.RAM_1.mem[512]);
      $display(" input buffer = %h", CPU.RAM_1.mem[513]);
      $display(" input buffer = %h", CPU.RAM_1.mem[514]);
      $display(" input buffer = %h", CPU.RAM_1.mem[515]);
      $display(" input buffer = %h", CPU.RAM_1.mem[516]);
      $display(" input buffer = %h", CPU.RAM_1.mem[517]);
      $display(" input buffer = %h", CPU.RAM_1.mem[518]);
      $display(" input buffer = %h", CPU.RAM_1.mem[519]);
      $display(" input buffer = %h", CPU.RAM_1.mem[520]);
      $display(" input buffer = %h", CPU.RAM_1.mem[521]);
      $display(" input buffer = %h", CPU.RAM_1.mem[522]);
      $display(" input buffer = %h", CPU.RAM_1.mem[523]);
      $display(" input buffer = %h", CPU.RAM_1.mem[524]);
      $display(" input buffer = %h", CPU.RAM_1.mem[525]);
      $display(" input buffer = %h", CPU.RAM_1.mem[526]);
      $display(" input buffer = %h", CPU.RAM_1.mem[527]);
      $display(" input buffer = %h", CPU.RAM_1.mem[528]);
      $display(" input buffer = %h", CPU.RAM_1.mem[529]);
      $display(" input buffer = %h", CPU.RAM_1.mem[530]);
      $display(" input buffer = %h", CPU.RAM_1.mem[531]);
      $display(" input buffer = %h", CPU.RAM_1.mem[532]);






      




        #1000 $finish();
      	
    end

endmodule
